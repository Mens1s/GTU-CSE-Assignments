module Or_32Bit(output [31:0] out, input [31:0] a, input[31:0] b);

    or o0(out[0], b[0], a[0]);
    or o1(out[1], b[1], a[1]);
    or o2(out[2], b[2], a[2]); 
    or o3(out[3], b[3], a[3]);
    or o4(out[4], b[4], a[4]);
    or o5(out[5], b[5], a[5]);
    or o6(out[6], b[6], a[6]);
    or o7(out[7], b[7], a[7]);
    or o8(out[8], b[8], a[8]);
    or o9(out[9], b[9], a[9]);
    or o10(out[10], b[10], a[10]);
    or o11(out[11], b[11], a[11]);
    or o12(out[12], b[12], a[12]);
    or o13(out[13], b[13], a[13]);
    or o14(out[14], b[14], a[14]);
    or o15(out[15], b[15], a[15]);
    or o16(out[16], b[16], a[16]);
    or o17(out[17], b[17], a[17]);
    or o18(out[18], b[18], a[18]);
    or o19(out[19], b[19], a[19]);
    or o20(out[20], b[20], a[20]);
    or o21(out[21], b[21], a[21]);
    or o22(out[22], b[22], a[22]);
    or o23(out[23], b[23], a[23]);
    or o24(out[24], b[24], a[24]);
    or o25(out[25], b[25], a[25]);
    or o26(out[26], b[26], a[26]);
    or o27(out[27], b[27], a[27]);
    or o28(out[28], b[28], a[28]);
    or o29(out[29], b[29], a[29]);
    or o30(out[30], b[30], a[30]);
    or o31(out[31], b[31], a[31]);

endmodule