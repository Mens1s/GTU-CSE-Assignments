module Nor_32Bit(output [31:0] out, input [31:0] a, input[31:0] b);

    nor no0(out[0], b[0], a[0]);
    nor no1(out[1], b[1], a[1]);
    nor no2(out[2], b[2], a[2]); 
    nor no3(out[3], b[3], a[3]);
    nor no4(out[4], b[4], a[4]);
    nor no5(out[5], b[5], a[5]);
    nor no6(out[6], b[6], a[6]);
    nor no7(out[7], b[7], a[7]);
    nor no8(out[8], b[8], a[8]);
    nor no9(out[9], b[9], a[9]);
    nor no10(out[10], b[10], a[10]);
    nor no11(out[11], b[11], a[11]);
    nor no12(out[12], b[12], a[12]);
    nor no13(out[13], b[13], a[13]);
    nor no14(out[14], b[14], a[14]);
    nor no15(out[15], b[15], a[15]);
    nor no16(out[16], b[16], a[16]);
    nor no17(out[17], b[17], a[17]);
    nor no18(out[18], b[18], a[18]);
    nor no19(out[19], b[19], a[19]);
    nor no20(out[20], b[20], a[20]);
    nor no21(out[21], b[21], a[21]);
    nor no22(out[22], b[22], a[22]);
    nor no23(out[23], b[23], a[23]);
    nor no24(out[24], b[24], a[24]);
    nor no25(out[25], b[25], a[25]);
    nor no26(out[26], b[26], a[26]);
    nor no27(out[27], b[27], a[27]);
    nor no28(out[28], b[28], a[28]);
    nor no29(out[29], b[29], a[29]);
    nor no30(out[30], b[30], a[30]);
    nor no31(out[31], b[31], a[31]);

endmodule