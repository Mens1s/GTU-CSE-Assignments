module OneBit_To_32Bit(
    output [31:0] result,
    input [0:0] wire1
);
    or or1(result[31], wire1[0], wire1[0]);
    or or2(result[30], wire1[0], wire1[0]);
    or or3(result[29], wire1[0], wire1[0]);
    or or4(result[28], wire1[0], wire1[0]);
    or or5(result[27], wire1[0], wire1[0]);
    or or6(result[26], wire1[0], wire1[0]);
    or or7(result[25], wire1[0], wire1[0]);
    or or8(result[24], wire1[0], wire1[0]);
    or or9(result[23], wire1[0], wire1[0]);
    or or10(result[22], wire1[0], wire1[0]);
    or or11(result[21], wire1[0], wire1[0]);
    or or12(result[20], wire1[0], wire1[0]);
    or or13(result[19], wire1[0], wire1[0]);
    or or14(result[18], wire1[0], wire1[0]);
    or or15(result[17], wire1[0], wire1[0]);
    or or16(result[16], wire1[0], wire1[0]);
    or or17(result[15], wire1[0], wire1[0]);
    or or18(result[14], wire1[0], wire1[0]);
    or or19(result[13], wire1[0], wire1[0]);
    or or20(result[12], wire1[0], wire1[0]);
    or or21(result[11], wire1[0], wire1[0]);
    or or22(result[10], wire1[0], wire1[0]);
    or or23(result[9], wire1[0], wire1[0]);
    or or24(result[8], wire1[0], wire1[0]);
    or or25(result[7], wire1[0], wire1[0]);
    or or26(result[6], wire1[0], wire1[0]);
    or or27(result[5], wire1[0], wire1[0]);
    or or28(result[4], wire1[0], wire1[0]);
    or or29(result[3], wire1[0], wire1[0]);
    or or30(result[2], wire1[0], wire1[0]);
    or or31(result[1], wire1[0], wire1[0]);
    or or32(result[0], wire1[0], wire1[0]);


endmodule