module And_32Bit (output [31:0] out, input [31:0] a, input [31:0] b);

    and a0(out[0], b[0], a[0]);
    and a1(out[1], b[1], a[1]);
    and a2(out[2], b[2], a[2]);
    and a3(out[3], b[3], a[3]);
    and a4(out[4], b[4], a[4]);
    and a5(out[5], b[5], a[5]);
    and a6(out[6], b[6], a[6]);
    and a7(out[7], b[7], a[7]);
    and a8(out[8], b[8], a[8]);
    and a9(out[9], b[9], a[9]);
    and a10(out[10], b[10], a[10]);
    and a11(out[11], b[11], a[11]);
    and a12(out[12], b[12], a[12]);
    and a13(out[13], b[13], a[13]);
    and a14(out[14], b[14], a[14]);
    and a15(out[15], b[15], a[15]);
    and a16(out[16], b[16], a[16]);
    and a17(out[17], b[17], a[17]);
    and a18(out[18], b[18], a[18]);
    and a19(out[19], b[19], a[19]);
    and a20(out[20], b[20], a[20]);
    and a21(out[21], b[21], a[21]);
    and a22(out[22], b[22], a[22]);
    and a23(out[23], b[23], a[23]);
    and a24(out[24], b[24], a[24]);
    and a25(out[25], b[25], a[25]);
    and a26(out[26], b[26], a[26]);
    and a27(out[27], b[27], a[27]);
    and a28(out[28], b[28], a[28]);
    and a29(out[29], b[29], a[29]);
    and a30(out[30], b[30], a[30]);
    and a31(out[31], b[31], a[31]);

endmodule